`timescale 1ps/1ps
module InstructionMemory(input [31:0]address,output reg[31:0] instruction);
  reg [7:0] IM[127:0];
	initial begin
	  IM[0] <= 8'b 00000000;
 		IM[1] <= 8'b 00000000;
 		IM[2] <= 8'b 00001000;
 		IM[3] <= 8'b 00100000;
 		IM[4] <= 8'b 00100000;
 		IM[5] <= 8'b 00100001;
 		IM[6] <= 8'b 00000011;
 		IM[7] <= 8'b 11101000;
 		IM[8] <= 8'b 00000000;
 		IM[9] <= 8'b 00000000;
 		IM[10] <= 8'b 00010000;
 		IM[11] <= 8'b 00100000;
 		IM[12] <= 8'b 00100000;
 		IM[13] <= 8'b 01000010;
 		IM[14] <= 8'b 00000100;
 		IM[15] <= 8'b 00010000;
		IM[16] <= 8'b 00000000;
		IM[17] <= 8'b 00000000;
		IM[18] <= 8'b 00011000;
		IM[19] <= 8'b 00100000;
		IM[20] <= 8'b 00010000;
		IM[21] <= 8'b 00100010;
		IM[22] <= 8'b 00000000;
		IM[23] <= 8'b 00000100;
		IM[24] <= 8'b 10001100;
		IM[25] <= 8'b 00100100;
		IM[26] <= 8'b 00000000;
		IM[27] <= 8'b 00000000;
		IM[28] <= 8'b 00000000;
		IM[29] <= 8'b 01100100;
		IM[30] <= 8'b 00011000;
		IM[31] <= 8'b 00100000;
		IM[32] <= 8'b 00100000;
		IM[33] <= 8'b 00100001;
		IM[34] <= 8'b 00000000;
		IM[35] <= 8'b 00000100;
		IM[36] <= 8'b 00001000;
		IM[37] <= 8'b 00000000;
		IM[38] <= 8'b 00000000;
		IM[39] <= 8'b 00000101;
//---------------------------------- 2 ----------------------------------------------
    
    //lui r8 ,1000......0
    {IM[40], IM[41], IM[42], IM[43]} <= {6'd15,5'd0,5'd8,16'b1000000000000000};
    //lw r2 1000 r0
		{IM[44], IM[45], IM[46], IM[47]} <= {6'd35,5'd0,5'd2,16'd1000};
		//addi r9,r0,0
		{IM[48], IM[49], IM[50], IM[51]} <= {6'd8,5'd0,5'd9,16'd0};
		//addi r6,r0,0
		{IM[52], IM[53], IM[54], IM[55]} <= {6'd8,5'd0,5'd6,16'd0};
		//addi r7,r0,20
		{IM[56], IM[57], IM[58], IM[59]} <= {6'd8,5'd0,5'd7,16'd20};
		//lw r1,1000,r6
		{IM[60], IM[61], IM[62], IM[63]} <= {6'd35,5'd6,5'd1,16'd1000};
		//sub r4,r2,r1
		{IM[64], IM[65], IM[66], IM[67]} <= {6'd0,5'd2,5'd1,5'd4,5'd0,6'd34};
		//and r5,r4,r8
		{IM[68], IM[69], IM[70], IM[71]} <= {6'd0,5'd4,5'd8,5'd5,5'd0,6'd36};
		//breq r5,r0,mosbat
		{IM[72], IM[73], IM[74], IM[75]} <= {6'd4,5'd5,5'd0,16'd2};
		//add r2,r0,r1
		{IM[76], IM[77], IM[78], IM[79]} <= {6'd0,5'd0,5'd1,5'd2,5'd0,6'd32};
		//add r3,r0,r9
		{IM[80], IM[81], IM[82], IM[83]} <= {6'd0,5'd0,5'd9,5'd3,5'd0,6'd32};
		//addi r9,r9,r1
		{IM[84], IM[85], IM[86], IM[87]} <= {6'd8,5'd9,5'd9,16'd1};
		//addi  r6,r6,4
		{IM[88], IM[89], IM[90], IM[91]} <= {6'd8,5'd6,5'd6,16'd4};
		//beq r9 r7 endfor
		{IM[92], IM[93], IM[94], IM[95]} <= {6'd4,5'd9,5'd7,16'd1};
		//jump for
		{IM[96], IM[97], IM[98], IM[99]} <= {6'd2,26'd15};
		//sw r2,2000(r0)
		{IM[100], IM[101], IM[102], IM[103]} <= {6'd43,5'd0,5'd2,16'd2000};
		//sw r3 2004(r0)
		{IM[104], IM[105], IM[106], IM[107]} <= {6'd43,5'd0,5'd3,16'd2004};


end
	always@(address)
		instruction = {IM[address], IM[address+1], IM[address+2], IM[address+3]};
endmodule